`timescale 1ns / 1ps
// Parameterized mux for a WISHBONE slave.
module wb_mux(
		sel_i,
		ack_i,
		rty_i,
		err_i,
		dat_i,
		dat_o
    );


endmodule
